package piso_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

//typedef uvm_config_db#(virtual piso_if) piso_vif_config;
`include "piso_item.sv"
`include "piso_monitor.sv"
`include "piso_sequencer.sv"
`include "piso_seq.sv"
`include "piso_driver.sv"
`include "piso_agent.sv"
`include "piso_sb.sv"
//`include "dummy_sb.sv"
`include "piso_env.sv"



endpackage
